
class pyhdl_object_type;

endclass
