
class pyhdl_uvm_type_info;

    /**
     */
    virtual function pyhdl_uvm_object create(uvm_object obj);
    endfunction

endclass
