
typedef class pyhdl_uvm_sequence_proxy_helper;
typedef class pyhdl_uvm_object_rgy;

class pyhdl_uvm_sequence_proxy #(
        type REQ=uvm_sequence_item, 
        type RSP=REQ, 
        type UserDataT=uvm_object,
        string PyClass="")
    extends uvm_sequence #(.REQ(REQ), .RSP(RSP));
    typedef pyhdl_uvm_sequence_proxy #(.REQ(REQ), .RSP(RSP), .PyClass(PyClass)) this_t;
    `uvm_object_param_utils(this_t);

    typedef pyhdl_uvm_sequence_proxy_helper #(.REQ(REQ), .RSP(RSP)) helper_t;

    string      pyclass = PyClass;
    UserDataT   userdata;
    helper_t    m_helper;

    function new(string name="pyhdl_uvm_sequence_proxy");
        super.new(name);
    endfunction

    virtual function uvm_object get_userdata();
        return userdata;
    endfunction

    task body();
        string modname, clsname;
        PyObject mod, cls;
        int i;

        // Ensure that the task scheduler is running
        pyhdl_if_start();

        if (pyclass == "") begin
            `uvm_fatal(get_name(), "No value specified for 'pyclass'");
        end

        for (i=pyclass.len()-1; i>=0; i--) begin
            if (pyclass[i] == ":") begin
                clsname = pyclass.substr(i+1, pyclass.len()-1);
                break;
            end
        end

        if (clsname == "") begin
            `uvm_fatal(get_name(), $sformatf("Failed to find '::' in pyclass %0s", pyclass))
        end

        for (; i>=0; i--) begin
            if (pyclass[i] != ":") begin
                break;
            end
        end

        modname = pyclass.substr(0, i);

        $display("modname=%0s clsname=%0s", modname, clsname);

        mod = PyImport_ImportModule(modname);
        if (mod == null) begin
            PyErr_Print();
            `uvm_fatal(get_name, $sformatf("Failed to load Python module %0s", modname));
            return;
        end

        cls = PyObject_GetAttrString(mod, clsname);

        if (cls == null) begin
            PyErr_Print();
            `uvm_fatal(get_name, $sformatf("Failed to find class %0s in Python module %0s", 
                clsname, modname));
            return;
        end

        m_helper = new(pyclass, cls);
        m_helper.m_proxy = this;
        m_helper.m_userdata = userdata;

        m_helper.body();
    endtask

endclass

class pyhdl_uvm_sequence_proxy_helper #(type REQ=uvm_sequence_item, type RSP=REQ)
        extends UvmSequenceProxy implements pyhdl_uvm_object_if;
    uvm_sequence_base       m_proxy;
    uvm_object              m_userdata;

    function new(string clsname, PyObject cls);
        PyObject impl_o, args;
        super.new();

        args = PyTuple_New(1);
        void'(PyTuple_SetItem(args, 0, m_obj));

        impl_o = PyObject_Call(cls, args, null);
        if (impl_o == null) begin
            PyErr_Print();
            $display("Fatal Error: Failed to construct user class %0s", clsname);
            $finish;
        end

        if (PyObject_SetAttrString(m_obj, "_impl", impl_o) != 0) begin
            PyErr_Print();
            $display("Fatal Error: Failed to set _impl on proxy wrapper");
            $finish;
        end
    endfunction

    virtual function uvm_object get_object();
        return m_proxy;
    endfunction

    virtual function string get_name();
        $display("get_name");
        return m_proxy.get_name();
    endfunction

    virtual function PyObject get_userdata();
        if (m_userdata != null) begin
            return pyhdl_uvm_object_rgy::inst().wrap(m_userdata);
        end else begin
            return None;
        end
    endfunction

    virtual function PyObject create_req();
        REQ req = REQ::type_id::create();
        return pyhdl_uvm_object_rgy::inst().wrap(req);
    endfunction

    virtual function PyObject create_rsp();
        RSP rsp = REQ::type_id::create();
        return pyhdl_uvm_object_rgy::inst().wrap(rsp);
    endfunction

    virtual task start_item(PyObject item);
        uvm_object item_o;
        uvm_sequence_item uvm_item;

        item_o = pyhdl_uvm_object_rgy::inst().get_object(item);
        if ($cast(uvm_item, item_o)) begin
            m_proxy.start_item(uvm_item);
        end else begin
            $display("Fatal: can't cast back to a sequence item");
        end
    endtask

    virtual task finish_item(PyObject item);
        uvm_object item_o;
        uvm_sequence_item uvm_item;

        item_o = pyhdl_uvm_object_rgy::inst().get_object(item);
        if ($cast(uvm_item, item_o)) begin
            m_proxy.finish_item(uvm_item);
        end else begin
            $display("Fatal: can't cast back to a sequence item");
        end
    endtask

endclass