
class vis_object_t;
endclass

