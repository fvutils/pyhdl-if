
typedef class vis_object_t;
class vis_component_t extends vis_object_t;

endclass
