`include "uvm_macros.svh"

module top;
  import uvm_pkg::*;
  import top_pkg::*;

  initial begin
    run_test();
  end

endmodule


