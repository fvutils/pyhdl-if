
module vpi_py_if_smoke;

initial begin
    $display("Hello World");
    $finish;
end

endmodule
