
class vis_component;

endclass

