/**
 * pyhdl_icall_api.sv
 *
 * Copyright 2024 Matthew Ballance and Contributors
 *
 * Licensed under the Apache License, Version 2.0 (the "License"); you may 
 * not use this file except in compliance with the License.  
 * You may obtain a copy of the License at:
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software 
 * distributed under the License is distributed on an "AS IS" BASIS, 
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  
 * See the License for the specific language governing permissions and 
 * limitations under the License.
 *
 * Created on:
 *     Author: 
 */
interface class ICallApi;

    pure virtual function PyObject invokeFunc(
        string              method,
        PyObject            args);

    pure virtual task invokeTask(
        output PyObject         retval,
        inout PyGILState_STATE  state,
        input string            method,
        input PyObject          args);

endclass