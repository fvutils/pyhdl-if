`include "uvm_macros.svh"

package pyhdl_if_uvm;
    import pyhdl_if::*;
    import uvm_pkg::*;


endpackage
