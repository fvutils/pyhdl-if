module top;
  import uvm_pkg::*;
  import reseed_pkg::*;

  initial begin
    run_test("reseed_test");
  end
endmodule
