
package pyhdl_if_vis;
    `include "vis_component.svh"
//         phase_listener pl = new("phase_listener");
endpackage
